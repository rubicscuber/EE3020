library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MovingLed_Basys3TB is
end entity MovingLed_Basys3TB;

--todo finnish this
architecture MovingLed_Basys3TB_ARCH of MovingLed_Basys3TB is
  
begin
  
  
  
end architecture MovingLed_Basys3TB_ARCH;
